import org.springframework.beans.factory.annotation.Autowired;
import org.springframework.stereotype.Service;
import java.util.List;

/**
 * Service层实现
 * 
 * @author XD.Wang
 * @date {new Date().format("yyyy-MM-dd")}
 */ 
@Service
public class {@cp}ServiceImpl implements {@cp}Service {

    @Autowired
    private {@cp}Mapper {@cl}Mapper;

    /**
     * 根据Example查询符合条件的结果列表
     * 
     * @param {@cl}Example 查询条件
     * @return 结果列表
     */
    @Override
    public List<{@cp}> select{@cp}ListByExample({@cp} {@cl}Example) {
        return {@cl}Mapper.select{@cp}ListByExample({@cl}Example);
    }

    /**
     * 根据DO参数查询符合条件的结果列表
     * 
     * @param {@cl} 查询条件
     * @return 结果列表
     */
    @Override
    public List<{@cp}> select{@cp}ListByParam({@cp} {@cl}) {
        return {@cl}Mapper.select{@cp}ListByParam({@cl});
    }

    /**
     * 根据ID查询符合条件的结果
     * 
     * @param id 主键
     * @return 结果
     */
    @Override
    public {@cp} select{@cp}ById(Long id) {
        return {@cl}Mapper.select{@cp}ById(id);
    }

    /**
     * 单条数据新增
     * 
     * @param {@cl} 待入库数据
     * @return 影响行数
     */
    @Override
    public Long insert{@cp}({@cp} {@cl}) {
        return {@cl}Mapper.insert{@cp}({@cl});
    }

    /**
     * 根据ID对单条数据更新
     * 
     * @param {@cl} 待入库数据
     * @return 影响行数
     */
    @Override
    public Long update{@cp}ById({@cp} {@cl}) {
        return {@cl}Mapper.update{@cp}ById({@cl});
    }

    /**
     * 根据主键删除
     * 
     * @param id 主键
     */
    @Override
    public void delete{@cp}ById(Long id) {
        {@cl}Mapper.delete{@cp}ById(id);
    }
    
}